module rand_num_rom(
	input clk,
	input [7:0] address,
	output reg [7:0] data
	);
	
	
	always @(posedge clk)
	begin
			case (address)
				8'd0 : data <= 8'd73;
				8'd1 : data <= 8'd95;
				8'd2 : data <= 8'd71;
				8'd3 : data <= 8'd127;
				8'd4 : data <= 8'd35;
				8'd5 : data <= 8'd21;
				8'd6 : data <= 8'd22;
				8'd7 : data <= 8'd17;
				8'd8 : data <= 8'd57;
				8'd9 : data <= 8'd63;
				8'd10 : data <= 8'd53;
				8'd11 : data <= 8'd99;
				8'd12 : data <= 8'd83;
				8'd13 : data <= 8'd100;
				8'd14 : data <= 8'd120;
				8'd15 : data <= 8'd124;
				8'd16 : data <= 8'd32;
				8'd17 : data <= 8'd26;
				8'd18 : data <= 8'd91;
				8'd19 : data <= 8'd21;
				8'd20 : data <= 8'd72;
				8'd21 : data <= 8'd116;
				8'd22 : data <= 8'd111;
				8'd23 : data <= 8'd67;
				8'd24 : data <= 8'd55;
				8'd25 : data <= 8'd89;
				8'd26 : data <= 8'd97;
				8'd27 : data <= 8'd71;
				8'd28 : data <= 8'd50;
				8'd29 : data <= 8'd140;
				8'd30 : data <= 8'd79;
				8'd31 : data <= 8'd139;
				8'd32 : data <= 8'd14;
				8'd33 : data <= 8'd98;
				8'd34 : data <= 8'd38;
				8'd35 : data <= 8'd62;
				8'd36 : data <= 8'd90;
				8'd37 : data <= 8'd145;
				8'd38 : data <= 8'd97;
				8'd39 : data <= 8'd56;
				8'd40 : data <= 8'd123;
				8'd41 : data <= 8'd92;
				8'd42 : data <= 8'd145;
				8'd43 : data <= 8'd100;
				8'd44 : data <= 8'd48;
				8'd45 : data <= 8'd126;
				8'd46 : data <= 8'd41;
				8'd47 : data <= 8'd33;
				8'd48 : data <= 8'd106;
				8'd49 : data <= 8'd60;
				8'd50 : data <= 8'd114;
				8'd51 : data <= 8'd55;
				8'd52 : data <= 8'd148;
				8'd53 : data <= 8'd56;
				8'd54 : data <= 8'd105;
				8'd55 : data <= 8'd98;
				8'd56 : data <= 8'd54;
				8'd57 : data <= 8'd35;
				8'd58 : data <= 8'd103;
				8'd59 : data <= 8'd122;
				8'd60 : data <= 8'd48;
				8'd61 : data <= 8'd89;
				8'd62 : data <= 8'd61;
				8'd63 : data <= 8'd108;
				8'd64 : data <= 8'd132;
				8'd65 : data <= 8'd30;
				8'd66 : data <= 8'd111;
				8'd67 : data <= 8'd126;
				8'd68 : data <= 8'd70;
				8'd69 : data <= 8'd114;
				8'd70 : data <= 8'd79;
				8'd71 : data <= 8'd28;
				8'd72 : data <= 8'd133;
				8'd73 : data <= 8'd57;
				8'd74 : data <= 8'd97;
				8'd75 : data <= 8'd106;
				8'd76 : data <= 8'd103;
				8'd77 : data <= 8'd47;
				8'd78 : data <= 8'd72;
				8'd79 : data <= 8'd20;
				8'd80 : data <= 8'd22;
				8'd81 : data <= 8'd115;
				8'd82 : data <= 8'd89;
				8'd83 : data <= 8'd68;
				8'd84 : data <= 8'd32;
				8'd85 : data <= 8'd68;
				8'd86 : data <= 8'd27;
				8'd87 : data <= 8'd16;
				8'd88 : data <= 8'd110;
				8'd89 : data <= 8'd75;
				8'd90 : data <= 8'd119;
				8'd91 : data <= 8'd91;
				8'd92 : data <= 8'd78;
				8'd93 : data <= 8'd146;
				8'd94 : data <= 8'd114;
				8'd95 : data <= 8'd126;
				8'd96 : data <= 8'd10;
				8'd97 : data <= 8'd112;
				8'd98 : data <= 8'd81;
				8'd99 : data <= 8'd126;
				8'd100 : data <= 8'd72;
				8'd101 : data <= 8'd66;
				8'd102 : data <= 8'd104;
				8'd103 : data <= 8'd37;
				8'd104 : data <= 8'd68;
				8'd105 : data <= 8'd115;
				8'd106 : data <= 8'd77;
				8'd107 : data <= 8'd109;
				8'd108 : data <= 8'd97;
				8'd109 : data <= 8'd79;
				8'd110 : data <= 8'd88;
				8'd112 : data <= 8'd20;
				8'd113 : data <= 8'd83;
				8'd114 : data <= 8'd88;
				8'd115 : data <= 8'd96;
				8'd116 : data <= 8'd114;
				8'd117 : data <= 8'd125;
				8'd118 : data <= 8'd100;
				8'd119 : data <= 8'd78;
				8'd120 : data <= 8'd119;
				8'd121 : data <= 8'd78;
				8'd122 : data <= 8'd12;
				8'd123 : data <= 8'd23;
				8'd124 : data <= 8'd111;
				8'd125 : data <= 8'd66;
				8'd126 : data <= 8'd109;
				8'd127 : data <= 8'd34;
				8'd128 : data <= 8'd74;
				8'd129 : data <= 8'd134;
				8'd130 : data <= 8'd13;
				8'd131 : data <= 8'd82;
				8'd132 : data <= 8'd52;
				8'd133 : data <= 8'd15;
				8'd134 : data <= 8'd67;
				8'd135 : data <= 8'd32;
				8'd136 : data <= 8'd24;
				8'd137 : data <= 8'd114;
				8'd138 : data <= 8'd27;
				8'd139 : data <= 8'd31;
				8'd140 : data <= 8'd14;
				8'd141 : data <= 8'd84;
				8'd142 : data <= 8'd43;
				8'd143 : data <= 8'd73;
				8'd144 : data <= 8'd91;
				
			endcase 
	
	end 
	
endmodule 